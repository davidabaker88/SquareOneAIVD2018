// nios_system.v

// Generated using ACDS version 17.0 602

`timescale 1 ps / 1 ps
module nios_system (
		input  wire [8:0]  blsensor_export,        //        blsensor.export
		input  wire [8:0]  brsensor_export,        //        brsensor.export
		input  wire [3:0]  challengeselect_export, // challengeselect.export
		input  wire        clk_clk,                //             clk.clk
		output wire [6:0]  drivespeed_export,      //      drivespeed.export
		input  wire [31:0] encoderincm_export,     //     encoderincm.export
		output wire        encoderreset_export,    //    encoderreset.export
		input  wire [8:0]  flsensor_export,        //        flsensor.export
		input  wire [8:0]  frsensor_export,        //        frsensor.export
		input  wire        greenlight_export,      //      greenlight.export
		output wire [7:0]  leds_export,            //            leds.export
		input  wire [8:0]  lsensor_export,         //         lsensor.export
		input  wire        redlight_export,        //        redlight.export
		input  wire        reset_reset_n,          //           reset.reset_n
		output wire        reverse_export,         //         reverse.export
		input  wire [8:0]  rsensor_export,         //         rsensor.export
		input  wire [7:0]  switches_export,        //        switches.export
		output wire [8:0]  targetdirection_export, // targetdirection.export
		input  wire        yellowlight_export      //     yellowlight.export
	);

	wire  [31:0] nios2_processor_data_master_readdata;                            // mm_interconnect_0:nios2_processor_data_master_readdata -> nios2_processor:d_readdata
	wire         nios2_processor_data_master_waitrequest;                         // mm_interconnect_0:nios2_processor_data_master_waitrequest -> nios2_processor:d_waitrequest
	wire         nios2_processor_data_master_debugaccess;                         // nios2_processor:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:nios2_processor_data_master_debugaccess
	wire  [18:0] nios2_processor_data_master_address;                             // nios2_processor:d_address -> mm_interconnect_0:nios2_processor_data_master_address
	wire   [3:0] nios2_processor_data_master_byteenable;                          // nios2_processor:d_byteenable -> mm_interconnect_0:nios2_processor_data_master_byteenable
	wire         nios2_processor_data_master_read;                                // nios2_processor:d_read -> mm_interconnect_0:nios2_processor_data_master_read
	wire         nios2_processor_data_master_write;                               // nios2_processor:d_write -> mm_interconnect_0:nios2_processor_data_master_write
	wire  [31:0] nios2_processor_data_master_writedata;                           // nios2_processor:d_writedata -> mm_interconnect_0:nios2_processor_data_master_writedata
	wire  [31:0] nios2_processor_instruction_master_readdata;                     // mm_interconnect_0:nios2_processor_instruction_master_readdata -> nios2_processor:i_readdata
	wire         nios2_processor_instruction_master_waitrequest;                  // mm_interconnect_0:nios2_processor_instruction_master_waitrequest -> nios2_processor:i_waitrequest
	wire  [18:0] nios2_processor_instruction_master_address;                      // nios2_processor:i_address -> mm_interconnect_0:nios2_processor_instruction_master_address
	wire         nios2_processor_instruction_master_read;                         // nios2_processor:i_read -> mm_interconnect_0:nios2_processor_instruction_master_read
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;        // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;          // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest;       // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;           // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;              // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;             // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;         // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire  [31:0] mm_interconnect_0_nios2_processor_jtag_debug_module_readdata;    // nios2_processor:jtag_debug_module_readdata -> mm_interconnect_0:nios2_processor_jtag_debug_module_readdata
	wire         mm_interconnect_0_nios2_processor_jtag_debug_module_waitrequest; // nios2_processor:jtag_debug_module_waitrequest -> mm_interconnect_0:nios2_processor_jtag_debug_module_waitrequest
	wire         mm_interconnect_0_nios2_processor_jtag_debug_module_debugaccess; // mm_interconnect_0:nios2_processor_jtag_debug_module_debugaccess -> nios2_processor:jtag_debug_module_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_processor_jtag_debug_module_address;     // mm_interconnect_0:nios2_processor_jtag_debug_module_address -> nios2_processor:jtag_debug_module_address
	wire         mm_interconnect_0_nios2_processor_jtag_debug_module_read;        // mm_interconnect_0:nios2_processor_jtag_debug_module_read -> nios2_processor:jtag_debug_module_read
	wire   [3:0] mm_interconnect_0_nios2_processor_jtag_debug_module_byteenable;  // mm_interconnect_0:nios2_processor_jtag_debug_module_byteenable -> nios2_processor:jtag_debug_module_byteenable
	wire         mm_interconnect_0_nios2_processor_jtag_debug_module_write;       // mm_interconnect_0:nios2_processor_jtag_debug_module_write -> nios2_processor:jtag_debug_module_write
	wire  [31:0] mm_interconnect_0_nios2_processor_jtag_debug_module_writedata;   // mm_interconnect_0:nios2_processor_jtag_debug_module_writedata -> nios2_processor:jtag_debug_module_writedata
	wire         mm_interconnect_0_onchip_memory_s1_chipselect;                   // mm_interconnect_0:onchip_memory_s1_chipselect -> onchip_memory:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory_s1_readdata;                     // onchip_memory:readdata -> mm_interconnect_0:onchip_memory_s1_readdata
	wire  [15:0] mm_interconnect_0_onchip_memory_s1_address;                      // mm_interconnect_0:onchip_memory_s1_address -> onchip_memory:address
	wire   [3:0] mm_interconnect_0_onchip_memory_s1_byteenable;                   // mm_interconnect_0:onchip_memory_s1_byteenable -> onchip_memory:byteenable
	wire         mm_interconnect_0_onchip_memory_s1_write;                        // mm_interconnect_0:onchip_memory_s1_write -> onchip_memory:write
	wire  [31:0] mm_interconnect_0_onchip_memory_s1_writedata;                    // mm_interconnect_0:onchip_memory_s1_writedata -> onchip_memory:writedata
	wire         mm_interconnect_0_onchip_memory_s1_clken;                        // mm_interconnect_0:onchip_memory_s1_clken -> onchip_memory:clken
	wire  [31:0] mm_interconnect_0_switches_s1_readdata;                          // switches:readdata -> mm_interconnect_0:switches_s1_readdata
	wire   [1:0] mm_interconnect_0_switches_s1_address;                           // mm_interconnect_0:switches_s1_address -> switches:address
	wire         mm_interconnect_0_leds_s1_chipselect;                            // mm_interconnect_0:LEDs_s1_chipselect -> LEDs:chipselect
	wire  [31:0] mm_interconnect_0_leds_s1_readdata;                              // LEDs:readdata -> mm_interconnect_0:LEDs_s1_readdata
	wire   [1:0] mm_interconnect_0_leds_s1_address;                               // mm_interconnect_0:LEDs_s1_address -> LEDs:address
	wire         mm_interconnect_0_leds_s1_write;                                 // mm_interconnect_0:LEDs_s1_write -> LEDs:write_n
	wire  [31:0] mm_interconnect_0_leds_s1_writedata;                             // mm_interconnect_0:LEDs_s1_writedata -> LEDs:writedata
	wire  [31:0] mm_interconnect_0_encoderincm_s1_readdata;                       // encoderInCM:readdata -> mm_interconnect_0:encoderInCM_s1_readdata
	wire   [1:0] mm_interconnect_0_encoderincm_s1_address;                        // mm_interconnect_0:encoderInCM_s1_address -> encoderInCM:address
	wire  [31:0] mm_interconnect_0_frsensor_s1_readdata;                          // FRSensor:readdata -> mm_interconnect_0:FRSensor_s1_readdata
	wire   [1:0] mm_interconnect_0_frsensor_s1_address;                           // mm_interconnect_0:FRSensor_s1_address -> FRSensor:address
	wire  [31:0] mm_interconnect_0_flsensor_s1_readdata;                          // FLSensor:readdata -> mm_interconnect_0:FLSensor_s1_readdata
	wire   [1:0] mm_interconnect_0_flsensor_s1_address;                           // mm_interconnect_0:FLSensor_s1_address -> FLSensor:address
	wire  [31:0] mm_interconnect_0_lsensor_s1_readdata;                           // LSensor:readdata -> mm_interconnect_0:LSensor_s1_readdata
	wire   [1:0] mm_interconnect_0_lsensor_s1_address;                            // mm_interconnect_0:LSensor_s1_address -> LSensor:address
	wire  [31:0] mm_interconnect_0_rsensor_s1_readdata;                           // RSensor:readdata -> mm_interconnect_0:RSensor_s1_readdata
	wire   [1:0] mm_interconnect_0_rsensor_s1_address;                            // mm_interconnect_0:RSensor_s1_address -> RSensor:address
	wire  [31:0] mm_interconnect_0_blsensor_s1_readdata;                          // BLSensor:readdata -> mm_interconnect_0:BLSensor_s1_readdata
	wire   [1:0] mm_interconnect_0_blsensor_s1_address;                           // mm_interconnect_0:BLSensor_s1_address -> BLSensor:address
	wire         mm_interconnect_0_drivespeed_s1_chipselect;                      // mm_interconnect_0:driveSpeed_s1_chipselect -> driveSpeed:chipselect
	wire  [31:0] mm_interconnect_0_drivespeed_s1_readdata;                        // driveSpeed:readdata -> mm_interconnect_0:driveSpeed_s1_readdata
	wire   [1:0] mm_interconnect_0_drivespeed_s1_address;                         // mm_interconnect_0:driveSpeed_s1_address -> driveSpeed:address
	wire         mm_interconnect_0_drivespeed_s1_write;                           // mm_interconnect_0:driveSpeed_s1_write -> driveSpeed:write_n
	wire  [31:0] mm_interconnect_0_drivespeed_s1_writedata;                       // mm_interconnect_0:driveSpeed_s1_writedata -> driveSpeed:writedata
	wire  [31:0] mm_interconnect_0_brsensor_s1_readdata;                          // BRSensor:readdata -> mm_interconnect_0:BRSensor_s1_readdata
	wire   [1:0] mm_interconnect_0_brsensor_s1_address;                           // mm_interconnect_0:BRSensor_s1_address -> BRSensor:address
	wire         mm_interconnect_0_targetdirection_s1_chipselect;                 // mm_interconnect_0:targetDirection_s1_chipselect -> targetDirection:chipselect
	wire  [31:0] mm_interconnect_0_targetdirection_s1_readdata;                   // targetDirection:readdata -> mm_interconnect_0:targetDirection_s1_readdata
	wire   [1:0] mm_interconnect_0_targetdirection_s1_address;                    // mm_interconnect_0:targetDirection_s1_address -> targetDirection:address
	wire         mm_interconnect_0_targetdirection_s1_write;                      // mm_interconnect_0:targetDirection_s1_write -> targetDirection:write_n
	wire  [31:0] mm_interconnect_0_targetdirection_s1_writedata;                  // mm_interconnect_0:targetDirection_s1_writedata -> targetDirection:writedata
	wire  [31:0] mm_interconnect_0_redlight_s1_readdata;                          // redlight:readdata -> mm_interconnect_0:redlight_s1_readdata
	wire   [1:0] mm_interconnect_0_redlight_s1_address;                           // mm_interconnect_0:redlight_s1_address -> redlight:address
	wire  [31:0] mm_interconnect_0_yellowlight_s1_readdata;                       // yellowlight:readdata -> mm_interconnect_0:yellowlight_s1_readdata
	wire   [1:0] mm_interconnect_0_yellowlight_s1_address;                        // mm_interconnect_0:yellowlight_s1_address -> yellowlight:address
	wire  [31:0] mm_interconnect_0_greenlight_s1_readdata;                        // greenlight:readdata -> mm_interconnect_0:greenlight_s1_readdata
	wire   [1:0] mm_interconnect_0_greenlight_s1_address;                         // mm_interconnect_0:greenlight_s1_address -> greenlight:address
	wire         mm_interconnect_0_reverse_s1_chipselect;                         // mm_interconnect_0:reverse_s1_chipselect -> reverse:chipselect
	wire  [31:0] mm_interconnect_0_reverse_s1_readdata;                           // reverse:readdata -> mm_interconnect_0:reverse_s1_readdata
	wire   [1:0] mm_interconnect_0_reverse_s1_address;                            // mm_interconnect_0:reverse_s1_address -> reverse:address
	wire         mm_interconnect_0_reverse_s1_write;                              // mm_interconnect_0:reverse_s1_write -> reverse:write_n
	wire  [31:0] mm_interconnect_0_reverse_s1_writedata;                          // mm_interconnect_0:reverse_s1_writedata -> reverse:writedata
	wire         mm_interconnect_0_encoderreset_s1_chipselect;                    // mm_interconnect_0:encoderreset_s1_chipselect -> encoderreset:chipselect
	wire  [31:0] mm_interconnect_0_encoderreset_s1_readdata;                      // encoderreset:readdata -> mm_interconnect_0:encoderreset_s1_readdata
	wire   [1:0] mm_interconnect_0_encoderreset_s1_address;                       // mm_interconnect_0:encoderreset_s1_address -> encoderreset:address
	wire         mm_interconnect_0_encoderreset_s1_write;                         // mm_interconnect_0:encoderreset_s1_write -> encoderreset:write_n
	wire  [31:0] mm_interconnect_0_encoderreset_s1_writedata;                     // mm_interconnect_0:encoderreset_s1_writedata -> encoderreset:writedata
	wire  [31:0] mm_interconnect_0_challengeselect_s1_readdata;                   // ChallengeSelect:readdata -> mm_interconnect_0:ChallengeSelect_s1_readdata
	wire   [1:0] mm_interconnect_0_challengeselect_s1_address;                    // mm_interconnect_0:ChallengeSelect_s1_address -> ChallengeSelect:address
	wire         irq_mapper_receiver0_irq;                                        // jtag_uart:av_irq -> irq_mapper:receiver0_irq
	wire  [31:0] nios2_processor_d_irq_irq;                                       // irq_mapper:sender_irq -> nios2_processor:d_irq
	wire         rst_controller_reset_out_reset;                                  // rst_controller:reset_out -> [BLSensor:reset_n, BRSensor:reset_n, ChallengeSelect:reset_n, FLSensor:reset_n, FRSensor:reset_n, LEDs:reset_n, LSensor:reset_n, RSensor:reset_n, driveSpeed:reset_n, encoderInCM:reset_n, encoderreset:reset_n, greenlight:reset_n, irq_mapper:reset, jtag_uart:rst_n, mm_interconnect_0:nios2_processor_reset_n_reset_bridge_in_reset_reset, nios2_processor:reset_n, onchip_memory:reset, redlight:reset_n, reverse:reset_n, rst_translator:in_reset, switches:reset_n, targetDirection:reset_n, yellowlight:reset_n]
	wire         rst_controller_reset_out_reset_req;                              // rst_controller:reset_req -> [nios2_processor:reset_req, onchip_memory:reset_req, rst_translator:reset_req_in]
	wire         nios2_processor_jtag_debug_module_reset_reset;                   // nios2_processor:jtag_debug_module_resetrequest -> rst_controller:reset_in1

	nios_system_BLSensor blsensor (
		.clk      (clk_clk),                                //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address  (mm_interconnect_0_blsensor_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_blsensor_s1_readdata), //                    .readdata
		.in_port  (blsensor_export)                         // external_connection.export
	);

	nios_system_BLSensor brsensor (
		.clk      (clk_clk),                                //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address  (mm_interconnect_0_brsensor_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_brsensor_s1_readdata), //                    .readdata
		.in_port  (brsensor_export)                         // external_connection.export
	);

	nios_system_ChallengeSelect challengeselect (
		.clk      (clk_clk),                                       //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),               //               reset.reset_n
		.address  (mm_interconnect_0_challengeselect_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_challengeselect_s1_readdata), //                    .readdata
		.in_port  (challengeselect_export)                         // external_connection.export
	);

	nios_system_BLSensor flsensor (
		.clk      (clk_clk),                                //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address  (mm_interconnect_0_flsensor_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_flsensor_s1_readdata), //                    .readdata
		.in_port  (flsensor_export)                         // external_connection.export
	);

	nios_system_BLSensor frsensor (
		.clk      (clk_clk),                                //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address  (mm_interconnect_0_frsensor_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_frsensor_s1_readdata), //                    .readdata
		.in_port  (frsensor_export)                         // external_connection.export
	);

	nios_system_LEDs leds (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_leds_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_leds_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_leds_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_leds_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_leds_s1_readdata),   //                    .readdata
		.out_port   (leds_export)                           // external_connection.export
	);

	nios_system_BLSensor lsensor (
		.clk      (clk_clk),                               //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address  (mm_interconnect_0_lsensor_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_lsensor_s1_readdata), //                    .readdata
		.in_port  (lsensor_export)                         // external_connection.export
	);

	nios_system_BLSensor rsensor (
		.clk      (clk_clk),                               //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address  (mm_interconnect_0_rsensor_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_rsensor_s1_readdata), //                    .readdata
		.in_port  (rsensor_export)                         // external_connection.export
	);

	nios_system_driveSpeed drivespeed (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_drivespeed_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_drivespeed_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_drivespeed_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_drivespeed_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_drivespeed_s1_readdata),   //                    .readdata
		.out_port   (drivespeed_export)                           // external_connection.export
	);

	nios_system_encoderInCM encoderincm (
		.clk      (clk_clk),                                   //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address  (mm_interconnect_0_encoderincm_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_encoderincm_s1_readdata), //                    .readdata
		.in_port  (encoderincm_export)                         // external_connection.export
	);

	nios_system_encoderreset encoderreset (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_encoderreset_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_encoderreset_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_encoderreset_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_encoderreset_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_encoderreset_s1_readdata),   //                    .readdata
		.out_port   (encoderreset_export)                           // external_connection.export
	);

	nios_system_greenlight greenlight (
		.clk      (clk_clk),                                  //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address  (mm_interconnect_0_greenlight_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_greenlight_s1_readdata), //                    .readdata
		.in_port  (greenlight_export)                         // external_connection.export
	);

	nios_system_jtag_uart jtag_uart (
		.clk            (clk_clk),                                                   //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                   //               irq.irq
	);

	nios_system_nios2_processor nios2_processor (
		.clk                                   (clk_clk),                                                         //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                                 //                   reset_n.reset_n
		.reset_req                             (rst_controller_reset_out_reset_req),                              //                          .reset_req
		.d_address                             (nios2_processor_data_master_address),                             //               data_master.address
		.d_byteenable                          (nios2_processor_data_master_byteenable),                          //                          .byteenable
		.d_read                                (nios2_processor_data_master_read),                                //                          .read
		.d_readdata                            (nios2_processor_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (nios2_processor_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (nios2_processor_data_master_write),                               //                          .write
		.d_writedata                           (nios2_processor_data_master_writedata),                           //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (nios2_processor_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (nios2_processor_instruction_master_address),                      //        instruction_master.address
		.i_read                                (nios2_processor_instruction_master_read),                         //                          .read
		.i_readdata                            (nios2_processor_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (nios2_processor_instruction_master_waitrequest),                  //                          .waitrequest
		.d_irq                                 (nios2_processor_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (nios2_processor_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_nios2_processor_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_nios2_processor_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_nios2_processor_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_nios2_processor_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_nios2_processor_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_nios2_processor_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_nios2_processor_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_nios2_processor_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                                 // custom_instruction_master.readra
	);

	nios_system_onchip_memory onchip_memory (
		.clk        (clk_clk),                                       //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),            //       .reset_req
		.freeze     (1'b0)                                           // (terminated)
	);

	nios_system_greenlight redlight (
		.clk      (clk_clk),                                //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address  (mm_interconnect_0_redlight_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_redlight_s1_readdata), //                    .readdata
		.in_port  (redlight_export)                         // external_connection.export
	);

	nios_system_encoderreset reverse (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_reverse_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_reverse_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_reverse_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_reverse_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_reverse_s1_readdata),   //                    .readdata
		.out_port   (reverse_export)                           // external_connection.export
	);

	nios_system_switches switches (
		.clk      (clk_clk),                                //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address  (mm_interconnect_0_switches_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_switches_s1_readdata), //                    .readdata
		.in_port  (switches_export)                         // external_connection.export
	);

	nios_system_targetDirection targetdirection (
		.clk        (clk_clk),                                         //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                 //               reset.reset_n
		.address    (mm_interconnect_0_targetdirection_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_targetdirection_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_targetdirection_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_targetdirection_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_targetdirection_s1_readdata),   //                    .readdata
		.out_port   (targetdirection_export)                           // external_connection.export
	);

	nios_system_greenlight yellowlight (
		.clk      (clk_clk),                                   //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address  (mm_interconnect_0_yellowlight_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_yellowlight_s1_readdata), //                    .readdata
		.in_port  (yellowlight_export)                         // external_connection.export
	);

	nios_system_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                       (clk_clk),                                                         //                                     clk_0_clk.clk
		.nios2_processor_reset_n_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                                  // nios2_processor_reset_n_reset_bridge_in_reset.reset
		.nios2_processor_data_master_address                 (nios2_processor_data_master_address),                             //                   nios2_processor_data_master.address
		.nios2_processor_data_master_waitrequest             (nios2_processor_data_master_waitrequest),                         //                                              .waitrequest
		.nios2_processor_data_master_byteenable              (nios2_processor_data_master_byteenable),                          //                                              .byteenable
		.nios2_processor_data_master_read                    (nios2_processor_data_master_read),                                //                                              .read
		.nios2_processor_data_master_readdata                (nios2_processor_data_master_readdata),                            //                                              .readdata
		.nios2_processor_data_master_write                   (nios2_processor_data_master_write),                               //                                              .write
		.nios2_processor_data_master_writedata               (nios2_processor_data_master_writedata),                           //                                              .writedata
		.nios2_processor_data_master_debugaccess             (nios2_processor_data_master_debugaccess),                         //                                              .debugaccess
		.nios2_processor_instruction_master_address          (nios2_processor_instruction_master_address),                      //            nios2_processor_instruction_master.address
		.nios2_processor_instruction_master_waitrequest      (nios2_processor_instruction_master_waitrequest),                  //                                              .waitrequest
		.nios2_processor_instruction_master_read             (nios2_processor_instruction_master_read),                         //                                              .read
		.nios2_processor_instruction_master_readdata         (nios2_processor_instruction_master_readdata),                     //                                              .readdata
		.BLSensor_s1_address                                 (mm_interconnect_0_blsensor_s1_address),                           //                                   BLSensor_s1.address
		.BLSensor_s1_readdata                                (mm_interconnect_0_blsensor_s1_readdata),                          //                                              .readdata
		.BRSensor_s1_address                                 (mm_interconnect_0_brsensor_s1_address),                           //                                   BRSensor_s1.address
		.BRSensor_s1_readdata                                (mm_interconnect_0_brsensor_s1_readdata),                          //                                              .readdata
		.ChallengeSelect_s1_address                          (mm_interconnect_0_challengeselect_s1_address),                    //                            ChallengeSelect_s1.address
		.ChallengeSelect_s1_readdata                         (mm_interconnect_0_challengeselect_s1_readdata),                   //                                              .readdata
		.driveSpeed_s1_address                               (mm_interconnect_0_drivespeed_s1_address),                         //                                 driveSpeed_s1.address
		.driveSpeed_s1_write                                 (mm_interconnect_0_drivespeed_s1_write),                           //                                              .write
		.driveSpeed_s1_readdata                              (mm_interconnect_0_drivespeed_s1_readdata),                        //                                              .readdata
		.driveSpeed_s1_writedata                             (mm_interconnect_0_drivespeed_s1_writedata),                       //                                              .writedata
		.driveSpeed_s1_chipselect                            (mm_interconnect_0_drivespeed_s1_chipselect),                      //                                              .chipselect
		.encoderInCM_s1_address                              (mm_interconnect_0_encoderincm_s1_address),                        //                                encoderInCM_s1.address
		.encoderInCM_s1_readdata                             (mm_interconnect_0_encoderincm_s1_readdata),                       //                                              .readdata
		.encoderreset_s1_address                             (mm_interconnect_0_encoderreset_s1_address),                       //                               encoderreset_s1.address
		.encoderreset_s1_write                               (mm_interconnect_0_encoderreset_s1_write),                         //                                              .write
		.encoderreset_s1_readdata                            (mm_interconnect_0_encoderreset_s1_readdata),                      //                                              .readdata
		.encoderreset_s1_writedata                           (mm_interconnect_0_encoderreset_s1_writedata),                     //                                              .writedata
		.encoderreset_s1_chipselect                          (mm_interconnect_0_encoderreset_s1_chipselect),                    //                                              .chipselect
		.FLSensor_s1_address                                 (mm_interconnect_0_flsensor_s1_address),                           //                                   FLSensor_s1.address
		.FLSensor_s1_readdata                                (mm_interconnect_0_flsensor_s1_readdata),                          //                                              .readdata
		.FRSensor_s1_address                                 (mm_interconnect_0_frsensor_s1_address),                           //                                   FRSensor_s1.address
		.FRSensor_s1_readdata                                (mm_interconnect_0_frsensor_s1_readdata),                          //                                              .readdata
		.greenlight_s1_address                               (mm_interconnect_0_greenlight_s1_address),                         //                                 greenlight_s1.address
		.greenlight_s1_readdata                              (mm_interconnect_0_greenlight_s1_readdata),                        //                                              .readdata
		.jtag_uart_avalon_jtag_slave_address                 (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),           //                   jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write                   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),             //                                              .write
		.jtag_uart_avalon_jtag_slave_read                    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),              //                                              .read
		.jtag_uart_avalon_jtag_slave_readdata                (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),          //                                              .readdata
		.jtag_uart_avalon_jtag_slave_writedata               (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),         //                                              .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest             (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest),       //                                              .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect              (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),        //                                              .chipselect
		.LEDs_s1_address                                     (mm_interconnect_0_leds_s1_address),                               //                                       LEDs_s1.address
		.LEDs_s1_write                                       (mm_interconnect_0_leds_s1_write),                                 //                                              .write
		.LEDs_s1_readdata                                    (mm_interconnect_0_leds_s1_readdata),                              //                                              .readdata
		.LEDs_s1_writedata                                   (mm_interconnect_0_leds_s1_writedata),                             //                                              .writedata
		.LEDs_s1_chipselect                                  (mm_interconnect_0_leds_s1_chipselect),                            //                                              .chipselect
		.LSensor_s1_address                                  (mm_interconnect_0_lsensor_s1_address),                            //                                    LSensor_s1.address
		.LSensor_s1_readdata                                 (mm_interconnect_0_lsensor_s1_readdata),                           //                                              .readdata
		.nios2_processor_jtag_debug_module_address           (mm_interconnect_0_nios2_processor_jtag_debug_module_address),     //             nios2_processor_jtag_debug_module.address
		.nios2_processor_jtag_debug_module_write             (mm_interconnect_0_nios2_processor_jtag_debug_module_write),       //                                              .write
		.nios2_processor_jtag_debug_module_read              (mm_interconnect_0_nios2_processor_jtag_debug_module_read),        //                                              .read
		.nios2_processor_jtag_debug_module_readdata          (mm_interconnect_0_nios2_processor_jtag_debug_module_readdata),    //                                              .readdata
		.nios2_processor_jtag_debug_module_writedata         (mm_interconnect_0_nios2_processor_jtag_debug_module_writedata),   //                                              .writedata
		.nios2_processor_jtag_debug_module_byteenable        (mm_interconnect_0_nios2_processor_jtag_debug_module_byteenable),  //                                              .byteenable
		.nios2_processor_jtag_debug_module_waitrequest       (mm_interconnect_0_nios2_processor_jtag_debug_module_waitrequest), //                                              .waitrequest
		.nios2_processor_jtag_debug_module_debugaccess       (mm_interconnect_0_nios2_processor_jtag_debug_module_debugaccess), //                                              .debugaccess
		.onchip_memory_s1_address                            (mm_interconnect_0_onchip_memory_s1_address),                      //                              onchip_memory_s1.address
		.onchip_memory_s1_write                              (mm_interconnect_0_onchip_memory_s1_write),                        //                                              .write
		.onchip_memory_s1_readdata                           (mm_interconnect_0_onchip_memory_s1_readdata),                     //                                              .readdata
		.onchip_memory_s1_writedata                          (mm_interconnect_0_onchip_memory_s1_writedata),                    //                                              .writedata
		.onchip_memory_s1_byteenable                         (mm_interconnect_0_onchip_memory_s1_byteenable),                   //                                              .byteenable
		.onchip_memory_s1_chipselect                         (mm_interconnect_0_onchip_memory_s1_chipselect),                   //                                              .chipselect
		.onchip_memory_s1_clken                              (mm_interconnect_0_onchip_memory_s1_clken),                        //                                              .clken
		.redlight_s1_address                                 (mm_interconnect_0_redlight_s1_address),                           //                                   redlight_s1.address
		.redlight_s1_readdata                                (mm_interconnect_0_redlight_s1_readdata),                          //                                              .readdata
		.reverse_s1_address                                  (mm_interconnect_0_reverse_s1_address),                            //                                    reverse_s1.address
		.reverse_s1_write                                    (mm_interconnect_0_reverse_s1_write),                              //                                              .write
		.reverse_s1_readdata                                 (mm_interconnect_0_reverse_s1_readdata),                           //                                              .readdata
		.reverse_s1_writedata                                (mm_interconnect_0_reverse_s1_writedata),                          //                                              .writedata
		.reverse_s1_chipselect                               (mm_interconnect_0_reverse_s1_chipselect),                         //                                              .chipselect
		.RSensor_s1_address                                  (mm_interconnect_0_rsensor_s1_address),                            //                                    RSensor_s1.address
		.RSensor_s1_readdata                                 (mm_interconnect_0_rsensor_s1_readdata),                           //                                              .readdata
		.switches_s1_address                                 (mm_interconnect_0_switches_s1_address),                           //                                   switches_s1.address
		.switches_s1_readdata                                (mm_interconnect_0_switches_s1_readdata),                          //                                              .readdata
		.targetDirection_s1_address                          (mm_interconnect_0_targetdirection_s1_address),                    //                            targetDirection_s1.address
		.targetDirection_s1_write                            (mm_interconnect_0_targetdirection_s1_write),                      //                                              .write
		.targetDirection_s1_readdata                         (mm_interconnect_0_targetdirection_s1_readdata),                   //                                              .readdata
		.targetDirection_s1_writedata                        (mm_interconnect_0_targetdirection_s1_writedata),                  //                                              .writedata
		.targetDirection_s1_chipselect                       (mm_interconnect_0_targetdirection_s1_chipselect),                 //                                              .chipselect
		.yellowlight_s1_address                              (mm_interconnect_0_yellowlight_s1_address),                        //                                yellowlight_s1.address
		.yellowlight_s1_readdata                             (mm_interconnect_0_yellowlight_s1_readdata)                        //                                              .readdata
	);

	nios_system_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.sender_irq    (nios2_processor_d_irq_irq)       //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                                // reset_in0.reset
		.reset_in1      (nios2_processor_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk            (clk_clk),                                       //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),                // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req),            //          .reset_req
		.reset_req_in0  (1'b0),                                          // (terminated)
		.reset_req_in1  (1'b0),                                          // (terminated)
		.reset_in2      (1'b0),                                          // (terminated)
		.reset_req_in2  (1'b0),                                          // (terminated)
		.reset_in3      (1'b0),                                          // (terminated)
		.reset_req_in3  (1'b0),                                          // (terminated)
		.reset_in4      (1'b0),                                          // (terminated)
		.reset_req_in4  (1'b0),                                          // (terminated)
		.reset_in5      (1'b0),                                          // (terminated)
		.reset_req_in5  (1'b0),                                          // (terminated)
		.reset_in6      (1'b0),                                          // (terminated)
		.reset_req_in6  (1'b0),                                          // (terminated)
		.reset_in7      (1'b0),                                          // (terminated)
		.reset_req_in7  (1'b0),                                          // (terminated)
		.reset_in8      (1'b0),                                          // (terminated)
		.reset_req_in8  (1'b0),                                          // (terminated)
		.reset_in9      (1'b0),                                          // (terminated)
		.reset_req_in9  (1'b0),                                          // (terminated)
		.reset_in10     (1'b0),                                          // (terminated)
		.reset_req_in10 (1'b0),                                          // (terminated)
		.reset_in11     (1'b0),                                          // (terminated)
		.reset_req_in11 (1'b0),                                          // (terminated)
		.reset_in12     (1'b0),                                          // (terminated)
		.reset_req_in12 (1'b0),                                          // (terminated)
		.reset_in13     (1'b0),                                          // (terminated)
		.reset_req_in13 (1'b0),                                          // (terminated)
		.reset_in14     (1'b0),                                          // (terminated)
		.reset_req_in14 (1'b0),                                          // (terminated)
		.reset_in15     (1'b0),                                          // (terminated)
		.reset_req_in15 (1'b0)                                           // (terminated)
	);

endmodule
