module SonicSensorNetwork (E1,T1,E2,T2,E3,T3,E4,T4,E5,T5,E6,T6,Dist1,Dist2,Dist3,Dist4,Dist5,Dist6,reset,CLOCK_50)
input wire CLOCK_50;
//echo
input wire E1;
input wire E2;
input wire E3;
input wire E4;
input wire E5;
input wire E6;
//trigger
output wire T1;
output wire T2;
output wire T3;
output wire T4;
output wire T5;
output wire T6;

wire TS1;
wire TS2;

assign T1 = TS1;
assign T3 = TS1;
assign T5 = TS1;
assign T2 = TS2;
assign T4 = TS2;
assign T6 = TS2;

SonicSensorTrig SST(
	.CLOCK_50(CLOCK_50),
	.reset(reset),
	.Tset1(TS1),
	.Tset2(TS2)
	);
//TS1
SonicSensor SS1(
	.CLOCK_50(CLOCK_50),
	.trigger(TS1),
	.echo(E1),
	.distanceCM(Dist1),
	.reset_n(~reset)
	);
SonicSensor SS3(
	.CLOCK_50(CLOCK_50),
	.trigger(TS1),
	.echo(E3),
	.distanceCM(Dist3),
	.reset_n(~reset)
	);
SonicSensor SS5(
	.CLOCK_50(CLOCK_50),
	.trigger(TS1),
	.echo(E5),
	.distanceCM(Dist5),
	.reset_n(~reset)
	);
//TS2
SonicSensor SS2(
	.CLOCK_50(CLOCK_50),
	.trigger(TS2),
	.echo(E2),
	.distanceCM(Dist2),
	.reset_n(~reset)
	);
SonicSensor SS4(
	.CLOCK_50(CLOCK_50),
	.trigger(TS4),
	.echo(E4),
	.distanceCM(Dist4),
	.reset_n(~reset)
	);
SonicSensor SS6(
	.CLOCK_50(CLOCK_50),
	.trigger(TS6),
	.echo(E6),
	.distanceCM(Dist6),
	.reset_n(~reset)
	);
	
endmodule
