// Implements a simple Nios II system for the DE-series board.
// Inputs: SW7¡0 are parallel port inputs to the Nios II system
// CLOCK_50 is the system clock
// KEY0 is the active-low system reset
// Outputs: LEDR7¡0 are parallel port outputs from the Nios II system
module ledTest (CLOCK_50, SW, KEY, LEDR);

input CLOCK_50;
input [7:0] SW;
input [0:0] KEY;
output [7:0] LEDR;

wire encReset;
wire reverse;
wire [8:0] targetDriection;
wire [6:0] driveSpeedPercentage;
wire [31:0] encoderInCM;
wire [8:0] RSesnorInCMl
wire [8:0] LSesnorInCM;
wire [8:0] BLSensorInCM;
wire [8:0] BRSensorInCM;
wire [8:0] LSensorInCM;
wire [8:0] FRSensorInCMdrive
wire [7:0] leftMagnetic;
wire [7:0] rightMagnetic;
wire reset
wire redLight;
wire greenLight;
wire yellowLight;


// Instantiate the Nios II system module generated by the Qsys tool:
nios_system NiosII (
.clk_clk(CLOCK_50),
.reset_reset_n(KEY),
.switches_export(SW),
.leds_export(LEDR));

	nios_system u0 (
		.blsensorincm_export         (BLSensorInCM),         //         blsensorincm.export
		.brsensorincm_export         (BRSensorInCM),         //         brsensorincm.export
		.clk_clk                     (CLOCK_50),                     //                  clk.clk
		.drivespeedpercentage_export (driveSpeedPercentage), // drivespeedpercentage.export
		.encoderincm_export          (encoderInCM),          //          encoderincm.export
		.flsensorincm_export         (FLSensorInCM),         //         flsensorincm.export
		.frsensorincm_export         (FRSensorInCM),         //         frsensorincm.export
		.leftmagnetic_export         (leftMagnetic),         //         leftmagnetic.export
		.lsensorincm_export          (LSensorInCM),          //          lsensorincm.export
		.reset_reset_n               (reset),               //                reset.reset_n
		.reverse_export              (reverse),              //              reverse.export
		.rightmagnetic_export        (rightMagnetic),        //        rightmagnetic.export
		.rsensorincm_export          (RSensorInCM),          //          rsensorincm.export
		.swiveldirection_export      (<connected-to-swiveldirection_export>),      //      swiveldirection.export
		.swiveldistacne_export       (<connected-to-swiveldistacne_export>),       //       swiveldistacne.export
		.targetdirection_export      (targetDirection),      //      targetdirection.export
		.encoderreset_export         (encReset)          //         encoderreset.export
	);
	
CustomLogic CL(

.encoderReset(encReset)
.targetDirection(targetDirection)
.driveSpeedPercentage(driveSpeedPercentage)
.reverse(reverse)
.encoderInCM(encoderInCM)
.RSensorInCM(RSensorInCM)
.LSensorInCM(LSensorInCM)
.FLSensorIncM(FLSensorInCM)
.FRSensorInCM(FRSensorInCM)
.BLSensorInCM(BLSensorInCM)
.BRSensorInCM(BRSensorInCM)
.leftMagnetic(leftMagnetic)
.rightMagnetic(rightMagnetic)
.redLight(redLight)
.yellowLight(yellowLight)
.greenLight(greenLight)
.reset(reset))

endmodule
