module SonicSensorNetwork (E1,T1,E2,T2,E3,T3,E4,T4,E5,T5,E6,T6,Dist1,Dist2,Dist3,Dist4,Dist5,Dist6,reset,CLOCK_50)

input wire E1;
input wire E2;
input wire E3;
input wire E4;
input wire E5;
input wire E6;
output wire T1;
output wire T2;
output wire T3;
output wire T4;
output wire T5;
output wire T6;
