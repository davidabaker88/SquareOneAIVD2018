// Implements a simple Nios II system for the DE-series board.
// Inputs: SW7¡0 are parallel port inputs to the Nios II system
// CLOCK_50 is the system clock
// KEY0 is the active-low system reset
// Outputs: LEDR7¡0 are parallel port outputs from the Nios II system
module ledTest (CLOCK_50, SW, KEY, LEDR, HEX0, HEX1, HEX2, HEX3, HEX4, HEX5,GPIO_0,GPIO_1);

input wire CLOCK_50;
input wire [7:0] SW;
input wire [3:0] KEY;
output wire [9:0] LEDR;
inout wire [39:0] GPIO_0;
inout wire [39:0] GPIO_1;

output wire [6:0] HEX0; 
output wire [6:0] HEX1;
output wire[6:0] HEX2; 
output wire[6:0] HEX3; 
output wire[6:0] HEX4; 
output wire[6:0] HEX5;  

wire [31:0] encoderInCM;
wire EncoderReset;
wire [8:0] FRSensorInCM;
wire [8:0] FLSensorInCM;
wire [8:0] LSensorInCM;
wire [8:0] RSensorInCM;
wire [8:0] BLSensorInCM;
wire [8:0] BRSensorInCM;
wire redLight;
wire yellowLight;
wire greenLight;
wire [6:0] driveSpeed;
wire reverse;
wire [7:0] targetDirection;
wire [3:0] challengeSelect;
reg temp;

assign redLight = 'b1;//GPIO_1[1];
assign yellowLight = 'b1;// GPIO_1[2];
assign greenLight = 'b1;// GPIO_1[3];
//assign GPIO_1[10] = CLOCK_50;
assign GPIO_1[11] = 'b0;


//assign LEDR[5] = CLOCK_50;


// Instantiate the Nios II system module generated by the Qsys tool:
nios_system NiosII (
.clk_clk(CLOCK_50),
.reset_reset_n(KEY[0]),
.switches_export(SW),
.leds_export(),
.encoderincm_export(encoderInCM),
.frsensor_export(FRSensorInCM),
.flsensor_export(FLSensorInCM),
.lsensor_export(LSensorInCM),
.rsensor_export(RSensorInCM),
.blsensor_export(BLSensorInCM),
.brsensor_export(BRSensorInCM),
.redlight_export(redLight),
.yellowlight_export(yellowLight),
.greenlight_export(greenLight),
//outputs
.drivespeed_export(driveSpeed),
.reverse_export(reverse),
.encoderreset_export(EncoderReset),
.targetdirection_export(targetDirection),
.challengeselect_export(challengeSelect));

CustomLogic CL(
.CLOCK_50(CLOCK_50),
.EncoderReset(EncoderReset),
.targetDirection(targetDirection),
.driveSpeedPercentage(driveSpeed),
.reverse(reverse),
.encoderInCM(encoderInCM),
.RSensorInCM(RSensorInCM),
.LSensorInCM(LSensorInCM),
.FLSensorInCM(FLSensorInCM),
.FRSensorInCM(FRSensorInCM),
.BLSensorInCM(BLSensorInCM),
.BRSensorInCM(BRSensorInCM),
.leftMagnetic(),
.rightMagnetic(),
.redLight(redLight),
.yellowLight(yellowLight),
.greenLight(greenLight),
.swivelDirection      (),      //      swiveldirection.export
.swivelDistance       (),
.HEX0(HEX0),
.HEX1(HEX1),
.HEX2(HEX2),
.HEX3(HEX3),
.HEX4(HEX4),
.HEX5(HEX5),
.LEDR(LEDR),
.SW(SW),
.KEY(~KEY),
.GPIO_0(GPIO_0),
.GPIO_1(GPIO_1),
.challengeSelect(challengeSelect));



	

endmodule 